`ifndef _my_include_vh_
`define _my_include_vh_

`define W 300
`define LOG_W 9
`define DATA_LENGTH  16
`endif
